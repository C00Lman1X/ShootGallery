    ����          Assembly-CSharp   	SaveUsers   _hit_bullet_minute_second_scene                    dB   3