    ����          Assembly-CSharp   
Menu+Value   hitbulletminutesecond                   �A