    ����          Assembly-CSharp   Menu+LoadScenes   	nameScene      1